NET clk LOC = "B8"; # Bank = 0, Signal name = MCLK

NET S_OUT[6] LOC = "L14"; # Bank = 1, Signal name = CA
NET S_OUT[5] LOC = "H12"; # Bank = 1, Signal name = CB
NET S_OUT[4] LOC = "N14"; # Bank = 1, Signal name = CC
NET S_OUT[3] LOC = "N11"; # Bank = 2, Signal name = CD
NET S_OUT[2] LOC = "P12"; # Bank = 2, Signal name = CE
NET S_OUT[1] LOC = "L13"; # Bank = 1, Signal name = CF
NET S_OUT[0] LOC = "M12"; # Bank = 1, Signal name = CG

NET sw[7] LOC = "N3";  # Bank = 2, Signal name = SW7
NET sw[6]  LOC = "E2";  # Bank = 3, Signal name = SW6
NET sw[5]  LOC = "F3";  # Bank = 3, Signal name = SW5
NET sw[4] LOC = "G3";  # Bank = 3, Signal name = SW4
NET sw[3]  LOC = "B4";  # Bank = 3, Signal name = SW3
NET sw[2]  LOC = "K3";  # Bank = 3, Signal name = SW2
NET sw[1]  LOC = "L3";  # Bank = 3, Signal name = SW1
NET sw[0]  LOC = "P11";  # Bank = 2, Signal name = SW0

NET AN_out[3] LOC = "K14"; # Bank = 1, Signal name = AN3
NET AN_out[2] LOC = "M13"; # Bank = 1, Signal name = AN2
NET AN_out[1] LOC = "J12"; # Bank = 1, Signal name = AN1
NET AN_out[0] LOC = "F12"; # Bank = 1, Signal name = AN0


NET button[3] LOC = "A7";  # Bank = 1, Signal name = BTN3
NET button[2] LOC = "M4";  # Bank = 0, Signal name = BTN2
NET button[1] LOC = "C11"; # Bank = 2, Signal name = BTN1
NET button[0] LOC = "G12"; # Bank = 0, Signal name = BTN0


